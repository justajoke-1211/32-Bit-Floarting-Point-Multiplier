module mux1b(in, out);
  input in;
  output out;
  assign out =(in) ? 1:0;
endmodule

  
