module mul(in1, in2, mul_e, out);
  input[22:0] in1, in2;
  input mul_e;
  output[47:0] out;
  
endmodule
